-- # Testbench pour l'unité LWR (Learning With Rounding)