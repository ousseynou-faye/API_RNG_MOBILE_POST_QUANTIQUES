-- # Interface Hash SHAKE pour le wrapper VHDL 